../../dds_test.srcs/sources_1/new/fifo.sv