../../dds_test.srcs/sim_1/new/axis_width_converter_test.sv