../../dds_test.srcs/sources_1/new/lfsr16.sv