../../dds_test.srcs/sources_1/new/sample_buffer.sv