../../dds_test.srcs/sources_1/new/banked_sample_buffer.sv