../../dds_test.srcs/sources_1/new/axis_width_converter.sv