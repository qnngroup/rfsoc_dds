../../dds_test.srcs/sim_1/new/sample_discriminator_test.sv