../../dds_test.srcs/sim_1/new/banked_sample_buffer_test.sv