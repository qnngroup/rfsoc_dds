../../dds_test.srcs/sources_1/new/timetagging_discriminating_buffer.sv