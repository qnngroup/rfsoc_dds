../../dds_test.srcs/sources_1/new/adc_axis_mux.sv