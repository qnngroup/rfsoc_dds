../dds_test.srcs/sources_1/new/axis.sv