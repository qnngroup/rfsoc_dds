../../dds_test.srcs/sim_1/new/sim_util_pkg.sv