../../dds_test.srcs/sim_1/new/dac_prescaler_test.sv