../../dds_test.srcs/sources_1/new/lmh6401_spi.sv