../../dds_test.srcs/sim_1/new/timetagging_discriminating_buffer_test.sv