../../dds_test.srcs/sim_1/new/fifo_test.sv