../../dds_test.srcs/sources_1/new/axis_x2.sv