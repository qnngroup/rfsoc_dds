../../dds_test.srcs/sources_1/new/noise_event_tracker.sv