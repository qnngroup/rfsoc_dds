../../dds_test.srcs/sim_1/new/sample_buffer_test.sv