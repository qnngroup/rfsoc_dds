../../dds_test.srcs/sim_1/new/axis_differentiator_test.sv