../../dds_test.srcs/sources_1/new/dac_prescaler.sv